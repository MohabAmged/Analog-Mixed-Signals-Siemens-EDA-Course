* Under Damped
R1 1 2 60
L1 2 3 0.04
C1 3 0 11.11u
Vsrc 1 0 1v

.end

Linear Circuit
R1 1 2 5000
V1 1 0 AC 1
C1 2 0 150n
.End

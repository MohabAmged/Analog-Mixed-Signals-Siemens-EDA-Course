*Lap Part 2

*Op Amp subcircuit
.SUBCKT opamp 1 2 3
* Connections / / /
            * / / /
            * / / /
            * / / Vin-
            * / Vin+
            * /
     *     output node

* First Stage of the op amp

* Differential Inputs

* +Ve Terminal Open Current Source (Topology Requirement to have atleaset 2 connections to a node )
Iopen 2 0 0A

* -Ve Terminal Open Current Source (Topology Requirement to have atleaset 2 connections to a node )
Iopen1 3 0 0A


* Define the Current controled Voltage source controlled by the Differntial inputs
Gin 0 4 2 3 10

* Defining The Passive elements to get the required specs 10000 Gain and ugf 10 MHz
R1 4 0 1000
*G*R1=10000
C1 4 0 159.155n
* R*C = 1.5915E-4
* G*R=1+jwRC @ UGF

* First stage Completed


*  2nd Stage of the op amp

* Ideal Output Buffer

* Define The Voltage Controlled Voltage Source  with output equal to the voltage across the Rc Components
Eout 1 0 4 0 1

.ends opamp

Xop1 out in+ in- opamp

*Vsrc src 0 AC 1v

*RF out in- 10k

*RF2 src in- 1k
Vsrc in+ 0 AC 1v

R in- 0 1

*.TF V(out) Vsrc

.AC DEC 20 1HZ 30MEGHZ

.PROBE


.end


* Under Damped used as function input Netlists 

R1 1 2 60
L1 2 3 0.04
C1 3 0 11.11u
Vsrc 1 0 AC 1
.AC DEC 10 1 10000
.end

*VCCS TEST
R1 1 0 1000
C1 1 0 159.15n
G1 0 1 2 0 10
E1 3 0 1 0 1
R3 3 0 1000
V1 2 0 AC 1
R2 2 0 1000
.AC DEC 100 1 10000
.PROBE
.end

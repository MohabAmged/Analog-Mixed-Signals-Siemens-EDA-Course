Linear Circuit
R1 1 2 5000
VSrc 1 0 AC 1
C1 2 0 150n
.AC DEC 100 1 10000
.PRINT AC V(1) V(2)

.PLOT AC V(1) V(2)



.End

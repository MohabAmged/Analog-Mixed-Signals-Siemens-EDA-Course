5T OTA

* Include external file that contains MOSFET Model
.INCLUDE ee214b_hspice.sp
** Circuit Description **

* power supply
VDD 7 0 DC 1.8
* input

* Add lines here to add the input (voltage)sources
Vin+ 4 0 1.2 AC 0.5
Vin- 3 0 1.2 AC -0.5
* circuit
* 5T OTA
M1 6 4 2 2 nch L=280n W=3.2u
M2 5 3 2 2 nch L=280n W=3.2u
M3 6 5 7 7 pch L=1.9u W=37.24u
M4 5 5 7 7 pch L=1.9u W=37.24u
M5 2 1 0 0 nch L=1u W=9.598u
CL 6 0 500f
* Current Mirror
M6 1 1 0 0 nch L=1u W=9.598u M=0.5
Iref 7 1 22.35u




** Analysis Requests **
.op
.ac dec 10 1 10e9

** Outputs Requests **
.PROBE

.END
